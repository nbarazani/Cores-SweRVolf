0000100B0000000B
800025370000002B
01C5062308000E13
01D5002301B00E93
01C5062300300E13
01C5042308700E13
0000059700050223
0005828306058593
03C000EF0000102B
001585930000002B
FE0296E300058283
000002DB0000102B
02000293020000EF
000012DB018000EF
0000006F010000EF
00958593800015B7
020FFF9301450F83
00550023FE0F8CE3
5265775300008067
6F53657375462B56
0A736B636F722043
2068636E61724220
2C7265746E756F63
2068636E61724220
6F43206E656B6154
203D207265746E75
0000000000000000
